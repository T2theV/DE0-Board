Library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY seven_seg_hex_nibble IS
PORT(	in_vect: IN STD_LOGIC_VECTOR(3 downto 0);
		out_vect: OUT STD_LOGIC_VECTOR(6 downto 0));
END ENTITY seven_seg_hex_nibble;

ARCHITECTURE muxes of seven_seg_hex_nibble IS
Begin
with in_vect select
	out_vect <= "1000000" when "0000",
					"1111001" when "0001",
					"0100100" when "0010",
					"0110000" when "0011",
					"0011001" when "0100",
					"0010010" when "0101",
					"0000010" when "0110",
					"1111000" when "0111",
					"0000000" when "1000",
					"0010000" when "1001",
					"0001000" when "1010",
					"0000011" when "1011",
					"0100111" when "1100",
					"0100001" when "1101",
					"0000110" when "1110",
					"0001110" when "1111",
					"0000000" when others;

end ARCHITECTURE muxes;