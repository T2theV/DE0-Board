--Library IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.NUMERIC_STD.ALL;
--
--ENTITY SIGNED_DISP IS
--PORT(number: IN STD_LOGIC_VECTOR(15 downto 0);
--		)